// Verilog HDL for gates, inv _functional

module inv (Y, A);
    output Y;
    input A;

not (Y, A);

endmodule
