// Verilog HDL for basic_gates, xor2 _functional

module xor2 (Y, A, B);
    output Y;
    input A;
    input B;

xor (Y, A, B);

endmodule
