// Global nets module 

`celldefine
module cds_globals;


supply1 vdd_;

supply0 gnd_;

supply1 vcc_;


endmodule
`endcelldefine
