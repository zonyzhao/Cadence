// Verilog HDL for basic_gates, xnor2 _functional

module xnor2 (Y, A, B);
    output Y;
    input A;
    input B;

xnor (Y, A, B);

endmodule
