// Verilog HDL for basic_gates, trinv0 _functional

module trinv0 (Y, A, _EN);
    output Y;
    input A;
    input _EN;

notif0 (Y, A, _EN);

endmodule
