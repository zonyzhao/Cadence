// Global nets module 

`celldefine
module cds_globals;


supply1 vcc_;

supply0 gnd_;

supply1 vdd_;


endmodule
`endcelldefine
