// Global nets module 

`celldefine
module cds_globals;


supply1 vdd_;

supply1 vcc_;

supply0 gnd_;


endmodule
`endcelldefine
