// Global nets module 

`celldefine
module cds_globals;


supply0 gnd_;

supply1 vdd_;

supply1 vcc_;

supply1 vddd_;


endmodule
`endcelldefine
